/*
    File name: pkg_config.sv
    Description: Testbench for register file.
    Author: Marko Gjorgjievski
    Date: 13.01.2025
*/

package pkg_config;
    localparam int DATA_WIDTH = 32;
    localparam int NUM_REGISTER = 32;
endpackage